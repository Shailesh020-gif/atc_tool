

module act_tb_top;

endmodule
